`timescale 1ns / 1ps

module uartInterface(
    );


endmodule
