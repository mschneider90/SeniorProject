`timescale 1ns / 1ps

//Supports up to 8 devices on a bi-directional bus

module BusController #(parameter ADDR_WIDTH = 16,
                       parameter DATA_WIDTH = 16)
                       ();
                       


endmodule
