`timescale 1ns / 1ps

module tb_impl_micron_controller(input clk50MHz,
                                 input button_1,
                                 input button_2);

micron_controller sram_ctrl



endmodule
