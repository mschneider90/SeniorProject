`timescale 1ns / 1ps

module ps2_controller(input clk,
                      input data
							 );

endmodule
