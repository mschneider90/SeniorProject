`timescale 1ns / 1ps

module tb_vga_module();

VGA_module();


endmodule
